-- If you got this far, you have learned the basics about working with Sigasi.
--
-- Congratulations!
--
-- TODO "Set up your own project"
-- You are now ready to go and set up a project for your own VHDL code.
-- Go to this webpage to lean how (you can hold CTRL and click on the link):
-- http://www.sigasi.com/app/project-setup
