------------------------------------------------------------------------
--
-- Copyright 1996 by IEEE. All rights reserved.
--
-- This source file is an essential part of IEEE Std 1076.2-1996, IEEE Standard 
-- VHDL Mathematical Packages. This source file may not be copied, sold, or 
-- included with software that is sold without written permission from the IEEE
-- Standards Department. This source file may be used to implement this standard 
-- and may be distributed in compiled form in any manner so long as the 
-- compiled form does not allow direct decompilation of the original source file.
-- This source file may be copied for individual use between licensed users. 
-- This source file is provided on an AS IS basis. The IEEE disclaims ANY 
-- WARRANTY EXPRESS OR IMPLIED INCLUDING ANY WARRANTY OF MERCHANTABILITY 
-- AND FITNESS FOR USE FOR A PARTICULAR PURPOSE. The user of the source 
-- file shall indemnify and hold IEEE harmless from any damages or liability 
-- arising out of the use thereof.
--
-- Title:       Standard VHDL Mathematical Packages (IEEE Std 1076.2-1996,
--              MATH_COMPLEX)
--
-- Library:     This package shall be compiled into a library
--              symbolically named IEEE.
--
-- Developers:  IEEE DASC VHDL Mathematical Packages Working Group
--
-- Purpose:     This package defines a standard for designers to use in
--              describing VHDL models that make use of common COMPLEX
--              constants and common COMPLEX mathematical functions and
--              operators.
--
-- Limitation:  The values generated by the functions in this package may
--              vary from platform to platform, and the precision of results
--              is only guaranteed to be the minimum required by IEEE Std 1076-
--              1993.
--
-- Notes:
--              No declarations or definitions shall be included in, or
--              excluded from, this package.
--              The "package declaration" defines the types, subtypes, and
--              declarations of MATH_COMPLEX.
--              The standard mathematical definition and conventional meaning
--              of the mathematical functions that are part of this standard
--              represent the formal semantics of the implementation of the
--              MATH_COMPLEX package declaration.  The purpose of the
--              MATH_COMPLEX package body is to provide a guideline for
--              implementations to verify their implementation of MATH_COMPLEX.
--              Tool developers may choose to implement the package body in
--              the most efficient manner available to them.
--
-- -----------------------------------------------------------------------------
-- Version    : 1.5
-- Date       : 24 July 1996
-- -----------------------------------------------------------------------------

use work.math_real.all;

package math_complex is
    constant CopyRightNotice: string
      := "Copyright 1996 IEEE. All rights reserved.";

    -- Type Definitions

    type complex is
        record
                re: real;        -- Real part
                im: real;        -- Imaginary part
        end record;

    subtype positive_real is real range 0.0 to real'high;

    subtype principal_value is real range -MATH_PI to MATH_PI;

    type complex_polar is
        record
                mag: positive_real;    -- Magnitude
                arg: principal_value;  -- Angle in radians; -MATH_PI is illegal
        end record;

    -- Constant Definitions

    constant  MATH_CBASE_1: complex := complex'(1.0, 0.0);
    constant  MATH_CBASE_J: complex := complex'(0.0, 1.0);
    constant  MATH_CZERO: complex := complex'(0.0, 0.0);


    --
    -- Overloaded equality and inequality operators for complex_polar
    -- (equality and inequality operators for complex are predefined)
    --

    --```
    -- Purpose:
    --         Returns `true` if `l` is equal to `r` and returns `false` otherwise
    -- Special values:
    --         `complex_polar'(0.0, x) = complex_polar'(0.0, y) returns true`
    --         regardless of the value of `x` and `y`.
    -- Domain:
    --         `l` in `complex_polar` and `l.arg /= -MATH_PI` and
    --         `r` in `complex_polar` and `r.arg /= -MATH_PI`
    -- Error conditions:
    --         Error if `l.arg = -MATH_PI`
    --         Error if `r.arg = -MATH_PI`
    -- Range:
    --         `"="(l,r)` is either `true` or `false`
    -- Notes:
    --         None
    --```
    function "=" ( l: in complex_polar;  r: in complex_polar ) return boolean;

    --```
    -- Purpose:
    --         returns true if l is not equal to r and returns false
    --         otherwise
    -- Special values:
    --         complex_polar'(0.0, x) /= complex_polar'(0.0, y) returns
    --         false regardless of the value of x and y.
    -- Domain:
    --         l in complex_polar and l.arg /= -MATH_PI
    --         r in complex_polar and r.arg /= -MATH_PI
    -- Error conditions:
    --         Error if l.arg = -MATH_PI
    --         Error if r.arg = -MATH_PI
    -- Range:
    --         "/="(l,r) is either true or false
    -- Notes:
    --         None
    --```
    function "/=" ( l: in complex_polar;  r: in complex_polar ) return boolean;

    -- Function Declarations

    --```
    -- Purpose:
    --         Returns complex number x + iy
    -- Special values:
    --         None
    -- Domain:
    --         x in real
    --         y in real
    -- Error conditions:
    --         None
    -- Range:
    --         cmplx(x,y) is mathematically unbounded
    -- Notes:
    --         None
    --```
    function cmplx(x: in real;  y: in real:= 0.0 ) return complex;

    --```
    -- Purpose:
    --         Returns principal value of angle X; X in radians
    -- Special values:
    --         None
    -- Domain:
    --         x in real
    -- Error conditions:
    --         None
    -- Range:
    --         -MATH_PI < get_principal_value(x) <= MATH_PI
    -- Notes:
    --         None
    --```
    function get_principal_value(x: in real ) return principal_value;

    --```
    -- Purpose:
    --         Returns principal value complex_polar of z
    -- Special values:
    --         complex_to_polar(math_czero) = complex_polar'(0.0, 0.0)
    --         complex_to_polar(z) = complex_polar'(abs(z.im),
    --                              sign(z.im)*MATH_PI_OVER_2) if z.re = 0.0
    -- Domain:
    --         z in complex
    -- Error conditions:
    --         None
    -- Range:
    --         result.mag >= 0.0
    --         -MATH_PI < result.arg <= MATH_PI
    -- Notes:
    --         None
    --```
    function complex_to_polar(z: in complex ) return complex_polar;

    --```
    -- Purpose:
    --         Returns complex value of z
    -- Special values:
    --         None
    -- Domain:
    --         z in complex_polar and z.arg /= -MATH_PI
    -- Error conditions:
    --         Error if z.arg = -MATH_PI
    -- Range:
    --         polar_to_complex(z) is mathematically unbounded
    -- Notes:
    --         None
    --```
    function polar_to_complex(z: in complex_polar ) return complex;

    --```
    -- Purpose:
    --         Returns absolute value (magnitude) of z
    -- Special values:
    --         None
    -- Domain:
    --         z in complex
    -- Error conditions:
    --         None
    -- Range:
    --         abs(z) is mathematically unbounded
    -- Notes:
    --         abs(z) = sqrt(z.re*z.re + z.im*z.im)
    --```
    function "abs"(z: in complex ) return positive_real;

    --```
    -- Purpose:
    --         Returns absolute value (magnitude) of z
    -- Special values:
    --         None
    -- Domain:
    --         z in complex_polar and z.arg /= -MATH_PI
    -- Error conditions:
    --         Error if z.arg = -MATH_PI
    -- Range:
    --         abs(z) >= 0.0
    -- Notes:
    --         abs(z) = z.mag
    --```
    function "abs"(z: in complex_polar ) return positive_real;

    --```
    -- Purpose:
    --         Returns argument (angle) in radians of the principal
    --         value of z
    -- Special values:
    --         arg(z) = 0.0 if z.re >= 0.0 and z.im = 0.0
    --         arg(z) = sign(z.im)*MATH_PI_OVER_2 if z.re = 0.0
    --         arg(z) = MATH_PI if z.re < 0.0        and z.im = 0.0
    -- Domain:
    --         z in complex
    -- Error conditions:
    --         None
    -- Range:
    --         -MATH_PI < arg(z) <= MATH_PI
    -- Notes:
    --         arg(z) = arctan(z.im, z.re)
    --```
    function arg(z: in complex ) return principal_value;

    --```
    -- Purpose:
    --         Returns argument (angle) in radians of the principal
    --         value of z
    -- Special values:
    --         None
    -- Domain:
    --         z in complex_polar and z.arg /= -MATH_PI
    -- Error conditions:
    --         Error if z.arg = -MATH_PI
    -- Range:
    --         -MATH_PI < arg(z) <= MATH_PI
    -- Notes:
    --         arg(z) = z.arg
    --```
    function arg(z: in complex_polar ) return principal_value;

    --```
    -- Purpose:
    --         Returns unary minus of z
    -- Special values:
    --         None
    -- Domain:
    --         z in complex
    -- Error conditions:
    --         None
    -- Range:
    --         "-"(z) is mathematically unbounded
    -- Notes:
    --         Returns -x -jy for z= x + jy
    --```
    function "-" (z: in complex ) return complex;

    --```
    -- Purpose:
    --         Returns principal value of unary minus of z
    -- Special values:
    --         "-"(z) = complex_polar'(z.mag, MATH_PI) if z.arg = 0.0
    -- Domain:
    --         z in complex_polar and z.arg /= -MATH_PI
    -- Error conditions:
    --         Error if z.arg = -MATH_PI
    -- Range:
    --         result.mag >= 0.0
    --         -MATH_PI < result.arg <= MATH_PI
    -- Notes:
    --         Returns complex_polar'(z.mag, z.arg - sign(z.arg)*MATH_PI) if
    --                z.arg /= 0.0
    --```
    function "-" (z: in complex_polar ) return complex_polar;

    --```
    -- Purpose:
    --         Returns complex conjugate of z
    -- Special values:
    --         None
    -- Domain:
    --         Z in complex
    -- Error conditions:
    --         None
    -- Range:
    --         conj(z) is mathematically unbounded
    -- Notes:
    --         Returns x -jy for z= x + jy
    --```
    function conj (z: in complex) return complex;

    --```
    -- Purpose:
    --         Returns principal value of complex conjugate of Z
    -- Special values:
    --         conj(z) = complex_polar'(z.mag, MATH_PI) if z.arg = MATH_PI
    -- Domain:
    --         z in complex_polar and z.arg /= -MATH_PI
    -- Error conditions:
    --         error if z.arg = -MATH_PI
    -- Range:
    --         result.mag >= 0.0
    --         -MATH_PI < result.arg <= MATH_PI
    -- Notes:
    --         Returns complex_polar'(z.mag, -z.arg) if z.arg /= MATH_PI
    --```
    function conj (z: in complex_polar) return complex_polar;

    --```
    -- Purpose:
    --         Returns square root of z with positive real part
    --         or, if the real part is zero, the one with nonnegative
    --         imaginary part
    -- Special values:
    --         sqrt(math_czero) = math_czero
    -- Domain:
    --         z in complex
    -- Error conditions:
    --         None
    -- Range:
    --         sqrt(z) is mathematically unbounded
    -- Notes:
    --         None
    --```
    function sqrt(z: in complex ) return complex;

    --```
    -- Purpose:
    --         Returns square root of z with positive real part
    --         or, if the real part is zero, the one with nonnegative
    --         imaginary part
    -- Special values:
    --         sqrt(z) = complex_polar'(0.0, 0.0) if z.mag = 0.0
    -- Domain:
    --         z in complex_polar and z.arg /= -MATH_PI
    -- Error conditions:
    --         Error if z.arg = -MATH_PI
    -- Range:
    --         result.mag >= 0.0
    --         -MATH_PI < result.arg <= MATH_PI
    -- Notes:
    --         None
    --```
    function sqrt(z: in complex_polar ) return complex_polar;

    --```
    -- Purpose:
    --         Returns exponential of z
    -- Special values:
    --         exp(math_czero) = math_cbase_1
    --         exp(z) = -math_cbase_1 if z.re = 0.0 and abs(z.im) = MATH_PI
    --         exp(z) = sign(z.im)*math_cbase_j if z.re = 0.0 and
    --                                          abs(z.im) =  MATH_PI_OVER_2
    -- Domain:
    --         z in complex
    -- Error conditions:
    --         None
    -- Range:
    --         exp(z) is mathematically unbounded
    -- Notes:
    --         None
    --```
    function exp(z: in complex ) return complex;

    --```
    -- Purpose:
    --         Returns principal value of exponential of z
    -- Special values:
    --         exp(z) = complex_polar'(1.0, 0.0) if z.mag =0.0 and
    --                                                        z.arg = 0.0
    --         exp(z) = complex_polar'(1.0, MATH_PI) if z.mag = MATH_PI and
    --                                        abs(z.arg) = MATH_PI_OVER_2
    --         exp(z) = complex_polar'(1.0, MATH_PI_OVER_2) if
    --                                        z.mag = MATH_PI_OVER_2 and
    --                                        z.arg = MATH_PI_OVER_2
    --         exp(z) = complex_polar'(1.0, -MATH_PI_OVER_2) if
    --                                        z.mag = MATH_PI_OVER_2 and
    --                                        z.arg = -MATH_PI_OVER_2
    -- Domain:
    --         z in complex_polar and z.arg /= -MATH_PI
    -- Error conditions:
    --         Error if z.arg = -MATH_PI
    -- Range:
    --         result.mag >= 0.0
    --         -MATH_PI < result.arg <= MATH_PI
    -- Notes:
    --         None
    --```
    function exp(z: in complex_polar ) return complex_polar;

    --```
    -- Purpose:
    --         Returns natural logarithm of z
    -- Special values:
    --         log(math_cbase_1) = math_czero
    --         log(-math_cbase_1) = complex'(0.0, MATH_PI)
    --         log(math_cbase_j) = complex'(0.0, MATH_PI_OVER_2)
    --         log(-math_cbase_j) = complex'(0.0, -MATH_PI_OVER_2)
    --         log(z) = math_cbase_1 if z = complex'(math_e, 0.0)
    -- Domain:
    --         z in complex and abs(z) /= 0.0
    -- Error conditions:
    --         Error if abs(z) = 0.0
    -- Range:
    --         log(z) is mathematically unbounded
    -- Notes:
    --         None
    --```
    function log(z: in complex ) return complex;

    --```
    -- Purpose:
    --         Returns logarithm base 2 of z
    -- Special values:
    --         log2(math_cbase_1) = math_czero
    --         log2(z) = math_cbase_1 if z = complex'(2.0, 0.0)
    -- Domain:
    --         z in complex and abs(z) /= 0.0
    -- Error conditions:
    --         error if abs(z) = 0.0
    -- Range:
    --         log2(z) is mathematically unbounded
    -- Notes:
    --         None
    --```
    function log2(z: in complex ) return complex;

    --```
    -- Purpose:
    --         Returns logarithm base 10 of z
    -- Special values:
    --         log10(math_cbase_1) = math_czero
    --         log10(z) = math_cbase_1 if z = complex'(10.0, 0.0)
    -- Domain:
    --         z in complex and abs(z) /= 0.0
    -- Error conditions:
    --         Error if abs(z) = 0.0
    -- Range:
    --         log10(z) is mathematically unbounded
    -- Notes:
    --         None
    --```
    function log10(z: in complex ) return complex;

    --```
    -- Purpose:
    --         Returns principal value of natural logarithm of z
    -- Special values:
    --         log(z) = complex_polar'(0.0, 0.0) if z.mag = 1.0 and
    --                                             z.arg = 0.0
    --         log(z) = complex_polar'(MATH_PI, MATH_PI_OVER_2) if
    --                              z.mag = 1.0 and z.arg = MATH_PI
    --         log(z) = complex_polar'(MATH_PI_OVER_2, MATH_PI_OVER_2) if
    --                              z.mag = 1.0 and  z.arg = MATH_PI_OVER_2
    --         log(z) = complex_polar'(MATH_PI_OVER_2, -MATH_PI_OVER_2) if
    --                              z.mag = 1.0 and  z.arg = -MATH_PI_OVER_2
    --         log(z) = complex_polar'(1.0, 0.0) if z.mag = math_e and
    --                                             z.arg = 0.0
    -- Domain:
    --         z in complex_polar and z.arg /= -MATH_PI
    --         z.mag /= 0.0
    -- Error conditions:
    --         Error if z.arg = -MATH_PI
    --         Error if z.mag = 0.0
    -- Range:
    --         result.mag >= 0.0
    --         -MATH_PI < result.arg <= MATH_PI
    -- Notes:
    --         None
    --```
    function log(z: in complex_polar ) return complex_polar;

    -- Purpose:
    --         Returns principal value of logarithm base 2 of z
    -- Special values:
    --         log2(z) = complex_polar'(0.0, 0.0) if z.mag = 1.0 and
    --                                              z.arg = 0.0
    --         log2(z) = complex_polar'(1.0, 0.0) if z.mag = 2.0 and
    --                                             z.arg = 0.0
    -- Domain:
    --         z in complex_polar and z.arg /= -MATH_PI
    --         z.mag /= 0.0
    -- Error conditions:
    --         Error if z.arg = -MATH_PI
    --         Error if z.mag = 0.0
    -- Range:
    --         result.mag >= 0.0
    --         -MATH_PI < result.arg <= MATH_PI
    -- Notes:
    --        None
    --```
    function log2(z: in complex_polar ) return complex_polar;

    --```
    -- Purpose:
    --         Returns principal value of logarithm base 10 of z
    -- Special values:
    --         log10(z) = complex_polar'(0.0, 0.0) if z.mag = 1.0 and
    --                                               z.arg = 0.0
    --         log10(z) = complex_polar'(1.0, 0.0) if z.mag = 10.0 and
    --                                               z.arg = 0.0
    -- Domain:
    --         z in complex_polar and z.arg /= -MATH_PI
    --         z.mag /= 0.0
    -- Error conditions:
    --         error if z.arg = -MATH_PI
    --         error if z.mag = 0.0
    -- Range:
    --         result.mag >= 0.0
    --         -MATH_PI < result.arg <= MATH_PI
    -- Notes:
    --         None
    --```
    function log10(z: in complex_polar ) return complex_polar;

    --```
    -- Purpose:
    --         Returns logarithm base base of z
    -- Special values:
    --         log(math_cbase_1, base) = math_czero
    --         log(z,base) = math_cbase_1 if z = complex'(base, 0.0)
    -- Domain:
    --         z in complex and abs(z) /= 0.0
    --         base > 0.0
    --         base /= 1.0
    -- Error conditions:
    --         error if abs(z) = 0.0
    --         error if base <= 0.0
    --         error if base = 1.0
    -- Range:
    --         log(z,base) is mathematically unbounded
    -- Notes:
    --         None
    --```
    function log(z: in complex; base: in real) return complex;

    --```
    -- Purpose:
    --         Returns principal value of logarithm base base of z
    -- Special values:
    --         log(z, base) = complex_polar'(0.0, 0.0) if z.mag = 1.0 and
    --                                                z.arg = 0.0
    --         log(z, base) = complex_polar'(1.0, 0.0) if z.mag = base and
    --                                                z.arg = 0.0
    -- Domain:
    --         z in complex_polar and z.arg /= -MATH_PI
    --         z.mag /= 0.0
    --         base > 0.0
    --         base /= 1.0
    -- Error conditions:
    --         Error if z.arg = -MATH_PI
    --         Error if z.mag = 0.0
    --         Error if base <= 0.0
    --         Error if base = 1.0
    -- Range:
    --         result.mag >= 0.0
    --         -MATH_PI < result.arg <= MATH_PI
    -- Notes:
    --         None
    --```
    function log(z: in complex_polar; base: in real ) return complex_polar;

    --```
    -- Purpose:
    --         Returns sine of z
    -- Special values:
    --         sin(math_czero) = math_czero
    --         sin(z) = math_czero if z = complex'(MATH_PI, 0.0)
    -- Domain:
    --         z in complex
    -- Error conditions:
    --         None
    -- Range:
    --         abs(sin(z)) <= sqrt(sin(z.re)*sin(z.re) +
    --                                         sinh(z.im)*sinh(z.im))
    -- Notes:
    --         None
    --```
    function sin (z : in complex ) return complex;

    --```
    -- Purpose:
    --         Returns principal value of sine of z
    -- Special values:
    --         sin(z) = complex_polar'(0.0, 0.0) if z.mag = 0.0 and
    --                                            z.arg = 0.0
    --         sin(z) = complex_polar'(0.0, 0.0) if z.mag = MATH_PI and
    --                                            z.arg = 0.0
    -- Domain:
    --         z in complex_polar and z.arg /= -MATH_PI
    -- Error conditions:
    --         Error if z.arg = -MATH_PI
    -- Range:
    --         result.mag >= 0.0
    --         -MATH_PI < result.arg <= MATH_PI
    -- Notes:
    --         None
    --```
    function sin (z : in complex_polar ) return complex_polar;

    --```
    -- Purpose:
    --         Returns cosine of z
    -- Special values:
    --         cos(z) = math_czero if z = complex'(MATH_PI_OVER_2, 0.0)
    --         cos(z) = math_czero if z = complex'(-MATH_PI_OVER_2, 0.0)
    -- Domain:
    --         z in complex
    -- Error conditions:
    --         None
    -- Range:
    --         abs(cos(z)) <= sqrt(cos(z.re)*cos(z.re) +
    --                                         sinh(z.im)*sinh(z.im))
    -- Notes:
    --         None
    --```
    function  cos (z : in complex ) return complex;

    --```
    -- Purpose:
    --         Returns principal value of cosine of z
    -- Special values:
    --         cos(z) = complex_polar'(0.0, 0.0) if z.mag = MATH_PI_OVER_2
    --                                               and z.arg = 0.0
    --         cos(z) = complex_polar'(0.0, 0.0) if z.mag = MATH_PI_OVER_2
    --                                               and z.arg = MATH_PI
    -- Domain:
    --         z in complex_polar and z.arg /= -MATH_PI
    -- Error conditions:
    --         error if z.arg = -MATH_PI
    -- Range:
    --         result.mag >= 0.0
    --         -MATH_PI < result.arg <= MATH_PI
    -- Notes:
    --         None
    --```
    function  cos (z : in complex_polar ) return complex_polar;

    --```
    -- Purpose:
    --         Returns hyperbolic sine of z
    -- Special values:
    --         sinh(math_czero) = math_czero
    --         sinh(z) = math_czero if z.re = 0.0 and z.im = MATH_PI
    --         sinh(z) = math_cbase_j if z.re = 0.0 and
    --                                               z.im = MATH_PI_OVER_2
    --         sinh(z) = -math_cbase_j if z.re = 0.0 and
    --                                               z.im = -MATH_PI_OVER_2
    -- Domain:
    --         z in complex
    -- Error conditions:
    --         None
    -- Range:
    --         abs(sinh(z)) <= sqrt(sinh(z.re)*sinh(z.re) +
    --                                         sin(z.im)*sin(z.im))
    -- Notes:
    --         None
    --```
    function sinh (z : in complex ) return complex;

    --```
    -- Purpose:
    --         Returns principal value of hyperbolic sine of z
    -- Special values:
    --         sinh(z) = complex_polar'(0.0, 0.0) if z.mag = 0.0 and
    --                                            z.arg = 0.0
    --         sinh(z) = complex_polar'(0.0, 0.0) if z.mag = MATH_PI and
    --                                            z.arg = MATH_PI_OVER_2
    --         sinh(z) = complex_polar'(1.0, MATH_PI_OVER_2) if z.mag =
    --                         MATH_PI_OVER_2 and z.arg = MATH_PI_OVER_2
    --         sinh(z) = complex_polar'(1.0, -MATH_PI_OVER_2) if z.mag =
    --                         MATH_PI_OVER_2 and z.arg = -MATH_PI_OVER_2
    -- Domain:
    --         z in complex_polar and z.arg /= -MATH_PI
    -- Error conditions:
    --         Error if z.arg = -MATH_PI
    -- Range:
    --         result.mag >= 0.0
    --         -MATH_PI < result.arg <= MATH_PI
    -- Notes:
    --         None
    --```
    function sinh (z : in complex_polar ) return complex_polar;

    --```
    -- Purpose:
    --         Returns hyperbolic cosine of z
    -- Special values:
    --         cosh(math_czero) = math_cbase_1
    --         cosh(z) = -math_cbase_1 if z.re = 0.0 and z.im = MATH_PI
    --         cosh(z) = math_czero if z.re = 0.0 and z.im = MATH_PI_OVER_2
    --         cosh(z) = math_czero if z.re = 0.0 and z.im = -MATH_PI_OVER_2
    -- Domain:
    --         z in complex
    -- Error conditions:
    --         None
    -- Range:
    --         abs(cosh(z)) <= sqrt(sinh(z.re)*sinh(z.re) +
    --                                         cos(z.im)*cos(z.im))
    -- Notes:
    --         None
    --```
    function cosh (z : in complex ) return complex;

    --```
    -- Purpose:
    --         Returns principal value of hyperbolic cosine of z
    -- Special values:
    --         cosh(z) = complex_polar'(1.0, 0.0) if z.mag = 0.0 and
    --                                            z.arg = 0.0
    --         cosh(z) = complex_polar'(1.0, MATH_PI) if z.mag = MATH_PI and
    --                                            z.arg = MATH_PI_OVER_2
    --         cosh(z) = complex_polar'(0.0, 0.0) if z.mag =
    --                        MATH_PI_OVER_2 and z.arg = MATH_PI_OVER_2
    --         cosh(z) = complex_polar'(0.0, 0.0) if z.mag =
    --                        MATH_PI_OVER_2 and z.arg = -MATH_PI_OVER_2
    -- Domain:
    --         z in complex_polar and z.arg /= -MATH_PI
    -- Error conditions:
    --         Error if z.arg = -MATH_PI
    -- Range:
    --         result.mag >= 0.0
    --         -MATH_PI < result.arg <= MATH_PI
    -- Notes:
    --         None
    --```
    function cosh (z : in complex_polar ) return complex_polar;

    --
    -- Arithmetic Operators
    --

    --```
    -- Purpose:
    --         Returns arithmetic addition of l and r
    -- Special values:
    --         None
    -- Domain:
    --         l in complex
    --         r in complex
    -- Error conditions:
    --         None
    -- Range:
    --         "+"(z) is mathematically unbounded
    -- Notes:
    --         None
    --```
    function "+" ( l: in complex;  r: in complex ) return complex;

    --```
    -- Purpose:
    --         Returns arithmetic addition of l and r
    -- Special values:
    --         None
    -- Domain:
    --         l in real
    --         r in complex
    -- Error conditions:
    --         None
    -- Range:
    --         "+"(z) is mathematically unbounded
    -- Notes:
    --         None
    --```
    function "+" ( l: in real;     r: in complex ) return complex;

    --```
    -- Purpose:
    --         Returns arithmetic addition of l and r
    -- Special values:
    --         None
    -- Domain:
    --         l in complex
    --         r in real
    -- Error conditions:
    --         None
    -- Range:
    --         "+"(z) is mathematically unbounded
    -- Notes:
    --         None
    --```
    function "+" ( l: in complex;  r: in real ) return complex;

    --```
    -- Purpose:
    --         Returns arithmetic addition of l and r
    -- Special values:
    --         None
    -- Domain:
    --         l in complex_polar and l.arg /= -MATH_PI
    --         r in complex_polar and r.arg /= -MATH_PI
    -- Error conditions:
    --         Error if l.arg = -MATH_PI
    --         Error if r.arg = -MATH_PI
    -- Range:
    --         result.mag >= 0.0
    --         -MATH_PI < result.arg <= MATH_PI
    -- Notes:
    --         None
    --```
    function "+" ( l: in complex_polar; r: in complex_polar) return complex_polar;

    --```
    -- Purpose:
    --         Returns arithmetic addition of l and r
    -- Special values:
    --         None
    -- Domain:
    --         l in real
    --         r in complex_polar and r.arg /= -MATH_PI
    -- Error conditions:
    --         Error if r.arg = -MATH_PI
    -- Range:
    --         result.mag >= 0.0
    --         -MATH_PI < result.arg <= MATH_PI
    -- Notes:
    --         None
    --```
    function "+" ( l: in real;  r: in complex_polar) return complex_polar;

    --```
    -- Purpose:
    --         Returns arithmetic addition of l and r
    -- Special values:
    --         None
    -- Domain:
    --         l in complex_polar and l.arg /= -MATH_PI
    --         r in real
    -- Error conditions:
    --         Error if l.arg = -MATH_PI
    -- Range:
    --         result.mag >= 0.0
    --         -MATH_PI < result.arg <= MATH_PI
    -- Notes:
    --         None
    --```
    function "+" ( l: in complex_polar;  r: in real) return complex_polar;

    --```
    -- Purpose:
    --         Returns arithmetic subtraction of l minus r
    -- Special values:
    --         None
    -- Domain:
    --         l in complex
    --         r in complex
    -- Error conditions:
    --         None
    -- Range:
    --         "-"(z) is mathematically unbounded
    -- Notes:
    --         None
    --```
    function "-" ( l: in complex;  r: in complex ) return complex;

    --```
    -- Purpose:
    --         Returns arithmetic subtraction of l minus r
    -- Special values:
    --         None
    -- Domain:
    --         l in real
    --         r in complex
    -- Error conditions:
    --         None
    -- Range:
    --         "-"(z) is mathematically unbounded
    -- Notes:
    --         None
    --```
    function "-" ( l: in real;     r: in complex ) return complex;

    --```
    -- Purpose:
    --         Returns arithmetic subtraction of l minus r
    -- Special values:
    --         None
    -- Domain:
    --         l in complex
    --         r in real
    -- Error conditions:
    --         None
    -- Range:
    --         "-"(z) is mathematically unbounded
    -- Notes:
    --         None
    --```
    function "-" ( l: in complex;  r: in real )    return complex;

    --```
    -- Purpose:
    --         Returns arithmetic subtraction of l minus r
    -- Special values:
    --         None
    -- Domain:
    --         l in complex_polar and l.arg /= -MATH_PI
    --         r in complex_polar and r.arg /= -MATH_PI
    -- Error conditions:
    --         Error if l.arg = -MATH_PI
    --         Error if r.arg = -MATH_PI
    -- Range:
    --         result.mag >= 0.0
    --         -MATH_PI < result.arg <= MATH_PI
    -- Notes:
    --         None
    --```
    function "-" ( l: in complex_polar; r: in complex_polar) return complex_polar;

    --```
    -- Purpose:
    --         Returns arithmetic subtraction of l minus r
    -- Special values:
    --         None
    -- Domain:
    --         l in real
    --         r in complex_polar and r.arg /= -MATH_PI
    -- Error conditions:
    --         Error if r.arg = -MATH_PI
    -- Range:
    --         result.mag >= 0.0
    --         -MATH_PI < result.arg <= MATH_PI
    -- Notes:
    --         None
    --```
    function "-" ( l: in real;  r: in complex_polar) return complex_polar;

    --```
    -- Purpose:
    --         Returns arithmetic subtraction of l minus r
    -- Special values:
    --         None
    -- Domain:
    --         l in complex_polar and l.arg /= -MATH_PI
    --         r in real
    -- Error conditions:
    --         Error if l.arg = -MATH_PI
    -- Range:
    --         result.mag >= 0.0
    --         -MATH_PI < result.arg <= MATH_PI
    -- Notes:
    --         None
    --```
    function "-" ( l: in complex_polar;  r: in real) return complex_polar;

    --```
    -- Purpose:
    --         Returns arithmetic multiplication of l and r
    -- Special values:
    --         None
    -- Domain:
    --         l in complex
    --         r in complex
    -- Error conditions:
    --         None
    -- Range:
    --         "*"(z) is mathematically unbounded
    -- Notes:
    --         None
    --```
    function "*" ( l: in complex;  r: in complex ) return complex;

    --```
    -- Purpose:
    --         Returns arithmetic multiplication of l and r
    -- Special values:
    --         None
    -- Domain:
    --         l in real
    --         r in complex
    -- Error conditions:
    --         None
    -- Range:
    --         "*"(z) is mathematically unbounded
    -- Notes:
    --         None
    --```
    function "*" ( l: in real;  r: in complex ) return complex;

    --```
    -- Purpose:
    --         Returns arithmetic multiplication of l and r
    -- Special values:
    --         None
    -- Domain:
    --         l in complex
    --         r in real
    -- Error conditions:
    --         None
    -- Range:
    --         "*"(z) is mathematically unbounded
    -- Notes:
    --         None
    --```
    function "*" ( l: in complex;  r: in real )  return complex;

    --```
    -- Purpose:
    --         Returns arithmetic multiplication of l and r
    -- Special values:
    --         None
    -- Domain:
    --         l in complex_polar and l.arg /= -MATH_PI
    --         r in complex_polar and r.arg /= -MATH_PI
    -- Error conditions:
    --         Error if l.arg = -MATH_PI
    --         error if r.arg = -MATH_PI
    -- Range:
    --         result.mag >= 0.0
    --         -MATH_PI < result.arg <= MATH_PI
    -- Notes:
    --         None
    --```
    function "*" ( l: in complex_polar; r: in complex_polar) return complex_polar;

    --```
    -- Purpose:
    --         Returns arithmetic multiplication of l and r
    -- Special values:
    --         None
    -- Domain:
    --         l in real
    --         r in complex_polar and r.arg /= -MATH_PI
    -- Error conditions:
    --         Error if r.arg = -MATH_PI
    -- Range:
    --         result.mag >= 0.0
    --         -MATH_PI < result.arg <= MATH_PI
    -- Notes:
    --         None
    --```
    function "*" ( l: in real;  r: in complex_polar) return complex_polar;

    --```
    -- Purpose:
    --         Returns arithmetic multiplication of l and r
    -- Special values:
    --         None
    -- Domain:
    --         l in complex_polar and l.arg /= -MATH_PI
    --         r in real
    -- Error conditions:
    --         Error if l.arg = -MATH_PI
    -- Range:
    --         result.mag >= 0.0
    --         -MATH_PI < result.arg <= MATH_PI
    -- Notes:
    --         None
    --```
    function "*" ( l: in complex_polar;  r: in real) return complex_polar;

    --```
    -- Purpose:
    --         Returns arithmetic division of l by r
    -- Special values:
    --         None
    -- Domain:
    --         l in complex
    --         r in complex and r /= math_czero
    -- Error conditions:
    --         Error if r = math_czero
    -- Range:
    --         "/"(z) is mathematically unbounded
    -- Notes:
    --         None
    --```
    function "/" ( l: in complex;  r: in complex ) return complex;

    --```
    -- Purpose:
    --         Returns arithmetic division of l by r
    -- Special values:
    --         None
    -- Domain:
    --         l in real
    --         r in complex and r /= math_czero
    -- Error conditions:
    --         Error if r = math_czero
    -- Range:
    --         "/"(z) is mathematically unbounded
    -- Notes:
    --         None
    --```
    function "/" ( l: in real;  r: in complex ) return complex;

    --```
    -- Purpose:
    --         Returns arithmetic division of l by r
    -- Special values:
    --         None
    -- Domain:
    --         l in complex
    --         r in real and r /= 0.0
    -- Error conditions:
    --         Error if r = 0.0
    -- Range:
    --         "/"(z) is mathematically unbounded
    -- Notes:
    --         None
    --```
    function "/" ( l: in complex;  r: in real ) return complex;

    --```
    -- Purpose:
    --         Returns arithmetic division of l by r
    -- Special values:
    --         None
    -- Domain:
    --         l in complex_polar and l.arg /= -MATH_PI
    --         r in complex_polar and r.arg /= -MATH_PI
    --         r.mag > 0.0
    -- Error conditions:
    --         Error if r.mag <= 0.0
    --         Error if l.arg = -MATH_PI
    --         Error if r.arg = -MATH_PI
    -- Range:
    --         result.mag >= 0.0
    --         -MATH_PI < result.arg <= MATH_PI
    -- Notes:
    --         None
    --```
    function "/" ( l: in complex_polar; r: in complex_polar) return complex_polar;

    --```
    -- Purpose:
    --         Returns arithmetic division of l by r
    -- Special values:
    --         None
    -- Domain:
    --         l in real
    --         r in complex_polar and r.arg /= -MATH_PI
    --         r.mag > 0.0
    -- Error conditions:
    --         Error if r.mag <= 0.0
    --         Error if r.arg = -MATH_PI
    -- Range:
    --         result.mag >= 0.0
    --         -MATH_PI < result.arg <= MATH_PI
    -- Notes:
    --         None
    --```
    function "/" ( l: in real;  r: in complex_polar) return complex_polar;

    --```
    -- Purpose:
    --         Returns arithmetic division of l by r
    -- Special values:
    --         None
    -- Domain:
    --         l in complex_polar and l.arg /= -MATH_PI
    --         r /= 0.0
    -- Error conditions:
    --         error if l.arg = -MATH_PI
    --         error if r = 0.0
    -- Range:
    --         result.mag >= 0.0
    --         -MATH_PI < result.arg <= MATH_PI
    -- Notes:
    --         None
    --```
    function "/" ( l: in complex_polar;  r: in real) return complex_polar;

end package math_complex;
